module dummy;
endmodule 
